library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package op_code is
    type opc is (s_and,s_eor,s_sub,s_rsb,s_add,s_adc,s_sbc,s_rsc,s_tst,s_teq,s_cmp,s_cmn,s_orr,s_mov,s_bic,s_mvn);
end package ;

package body op_code is
    
end op_code;